{"bisBaseClass":"SpatialViewDefinition","viewDefinitionProps":{"classFullName":"BisCore:SpatialViewDefinition","id":"0x40000000060","jsonProperties":{"viewDetails":{"gridOrient":4,"gridPerRef":100,"gridSpaceX":0.1}},"code":{"spec":"0x1c","scope":"0x40000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x40000000007","categorySelectorId":"0x40000000063","displayStyleId":"0x40000000062","isPrivate":false,"description":"","cameraOn":true,"origin":[-34.29876483299998,34.72276642647075,-20.762995661518858],"extents":[109.9796056733849,51.11373077427796,129.45606652680968],"angles":{"pitch":-42.38875364730823,"roll":-55.48084033403707,"yaw":24.875625209910112},"camera":{"lens":45.87079213591108,"focusDist":129.95506652680584,"eye":[-77.12275597351177,-78.01360530134251,56.84001513058834]},"modelSelectorId":"0x40000000061"},"categorySelectorProps":{"classFullName":"BisCore:CategorySelector","id":"0x40000000063","code":{"spec":"0x8","scope":"0x40000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x40000000007","categories":["0x40000000008","0x4000000003f","0x40000000041","0x40000000043","0x40000000045","0x40000000047","0x40000000049","0x4000000004b","0x4000000004d","0x4000000004f","0x40000000051","0x40000000053","0x40000000055","0x40000000057","0x40000000059","0x4000000005b"]},"displayStyleProps":{"classFullName":"BisCore:DisplayStyle3d","id":"0x40000000062","jsonProperties":{"styles":{"hline":{"visible":{"ovrColor":true,"color":0,"pattern":0,"width":1},"hidden":{"ovrColor":true,"color":0,"pattern":3435973836,"width":1},"transThreshold":0.3},"sceneLights":{"ambient":{"intensity":20,"type":2},"sun":{"intensity":99415.46481844832,"type":1},"sunDir":[-6.123233995736766e-17,-3.749399456654644e-33,-1],"portrait":{"intensity":100,"intensity2":100,"type":4},"fstop":0.8570573925971985},"viewflags":{"grid":true,"noSolarLight":true,"noSourceLights":true,"renderMode":6,"visEdges":true},"environment":{"ground":{"aboveColor":32768,"belowColor":1262987,"display":false,"elevation":-0.01},"sky":{"display":false,"groundColor":8228728,"groundExponent":4,"image":{"texture":"0","type":0},"nadirColor":3880,"skyColor":16764303,"skyExponent":4,"zenithColor":16741686}}}},"code":{"spec":"0xa","scope":"0x40000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x40000000007"},"modelSelectorProps":{"classFullName":"BisCore:ModelSelector","id":"0x40000000061","code":{"spec":"0x11","scope":"0x40000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x40000000007","models":["0x40000000030"]}}