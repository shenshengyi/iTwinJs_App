{"bisBaseClass":"SpatialViewDefinition","viewDefinitionProps":{"classFullName":"BisCore:SpatialViewDefinition","id":"0x40000000060","jsonProperties":{"viewDetails":{"gridOrient":4,"gridPerRef":100,"gridSpaceX":0.1}},"code":{"spec":"0x1c","scope":"0x40000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x40000000007","categorySelectorId":"0x40000000063","displayStyleId":"0x40000000062","isPrivate":false,"description":"","cameraOn":true,"origin":[-47.885958497069964,18.03998925997445,-23.013418081201113],"extents":[106.24577326685984,49.378408091360065,125.54306272102079],"angles":{"pitch":-42.38875364730819,"roll":-55.48084033403707,"yaw":24.87562520991013},"camera":{"lens":45.87079213591113,"focusDist":125.54306272101888,"eye":[-89.59249292756566,-91.17264410557317,52.16382076096789]},"modelSelectorId":"0x40000000061"},"categorySelectorProps":{"classFullName":"BisCore:CategorySelector","id":"0x40000000063","code":{"spec":"0x8","scope":"0x40000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x40000000007","categories":["0x40000000008","0x4000000003f","0x40000000041","0x40000000043","0x40000000045","0x40000000047","0x40000000049","0x4000000004b","0x4000000004d","0x4000000004f","0x40000000051","0x40000000053","0x40000000055","0x40000000057","0x40000000059","0x4000000005b"]},"displayStyleProps":{"classFullName":"BisCore:DisplayStyle3d","id":"0x40000000062","jsonProperties":{"styles":{"hline":{"visible":{"ovrColor":true,"color":0,"pattern":0,"width":1},"hidden":{"ovrColor":true,"color":0,"pattern":3435973836,"width":1},"transThreshold":0.3},"sceneLights":{"ambient":{"intensity":20,"type":2},"sun":{"intensity":99415.46481844832,"type":1},"sunDir":[-6.123233995736766e-17,-3.749399456654644e-33,-1],"portrait":{"intensity":100,"intensity2":100,"type":4},"fstop":0.8570573925971985},"viewflags":{"grid":true,"noSolarLight":true,"noSourceLights":true,"renderMode":6,"visEdges":true},"environment":{"ground":{"aboveColor":32768,"belowColor":1262987,"display":false,"elevation":-0.01},"sky":{"display":false,"groundColor":8228728,"groundExponent":4,"image":{"texture":"0","type":0},"nadirColor":3880,"skyColor":16764303,"skyExponent":4,"zenithColor":16741686}}}},"code":{"spec":"0xa","scope":"0x40000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x40000000007"},"modelSelectorProps":{"classFullName":"BisCore:ModelSelector","id":"0x40000000061","code":{"spec":"0x11","scope":"0x40000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x40000000007","models":["0x40000000030"]}}