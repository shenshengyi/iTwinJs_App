{"bisBaseClass":"SpatialViewDefinition","viewDefinitionProps":{"classFullName":"BisCore:SpatialViewDefinition","id":"0x50000000060","jsonProperties":{"viewDetails":{"gridOrient":4,"gridPerRef":100,"gridSpaceX":0.1}},"code":{"spec":"0x1c","scope":"0x50000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x50000000007","categorySelectorId":"0x50000000063","displayStyleId":"0x50000000062","isPrivate":false,"description":"","cameraOn":true,"origin":[-47.07306090941197,25.473531897182443,-20.99484072670538],"extents":[101.06002004412802,46.96829584858903,118.91642750242274],"angles":{"pitch":-42.38875364730822,"roll":-55.48084033403712,"yaw":24.875625209910112},"camera":{"lens":45.87079213591103,"focusDist":119.41542750242158,"eye":[-86.42398774476716,-78.11972382297182,50.31443076374244]},"modelSelectorId":"0x50000000061"},"categorySelectorProps":{"classFullName":"BisCore:CategorySelector","id":"0x50000000063","code":{"spec":"0x8","scope":"0x50000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x50000000007","categories":["0x50000000008","0x5000000003f","0x50000000041","0x50000000043","0x50000000045","0x50000000047","0x50000000049","0x5000000004b","0x5000000004d","0x5000000004f","0x50000000051","0x50000000053","0x50000000055","0x50000000057","0x50000000059","0x5000000005b"]},"displayStyleProps":{"classFullName":"BisCore:DisplayStyle3d","id":"0x50000000062","jsonProperties":{"styles":{"hline":{"visible":{"ovrColor":true,"color":0,"pattern":0,"width":1},"hidden":{"ovrColor":true,"color":0,"pattern":3435973836,"width":1},"transThreshold":0.3},"sceneLights":{"ambient":{"intensity":20,"type":2},"sun":{"intensity":99415.46481844832,"type":1},"sunDir":[-6.123233995736766e-17,-3.749399456654644e-33,-1],"portrait":{"intensity":100,"intensity2":100,"type":4},"fstop":0.8570573925971985},"viewflags":{"grid":true,"noSolarLight":true,"noSourceLights":true,"renderMode":6,"visEdges":true},"environment":{"ground":{"aboveColor":32768,"belowColor":1262987,"display":false,"elevation":-0.01},"sky":{"display":false,"groundColor":8228728,"groundExponent":4,"image":{"texture":"0","type":0},"nadirColor":3880,"skyColor":16764303,"skyExponent":4,"zenithColor":16741686}}}},"code":{"spec":"0xa","scope":"0x50000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x50000000007"},"modelSelectorProps":{"classFullName":"BisCore:ModelSelector","id":"0x50000000061","code":{"spec":"0x11","scope":"0x50000000007","value":"3D Metric Design Model Views - View 1"},"model":"0x50000000007","models":["0x50000000030"]}}